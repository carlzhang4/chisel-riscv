module Regfile(
  input         clock,
  input         reset,
  input  [4:0]  io_w_addr,
  input  [31:0] io_w_data,
  input         io_w_en,
  input  [4:0]  io_r1_addr,
  output [31:0] io_r1_data,
  input         io_r1_en,
  input  [4:0]  io_r2_addr,
  output [31:0] io_r2_data,
  input         io_r2_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] registers_0; // @[Reg_file.scala 20:28]
  reg [31:0] registers_1; // @[Reg_file.scala 20:28]
  reg [31:0] registers_2; // @[Reg_file.scala 20:28]
  reg [31:0] registers_3; // @[Reg_file.scala 20:28]
  reg [31:0] registers_4; // @[Reg_file.scala 20:28]
  reg [31:0] registers_5; // @[Reg_file.scala 20:28]
  reg [31:0] registers_6; // @[Reg_file.scala 20:28]
  reg [31:0] registers_7; // @[Reg_file.scala 20:28]
  reg [31:0] registers_8; // @[Reg_file.scala 20:28]
  reg [31:0] registers_9; // @[Reg_file.scala 20:28]
  reg [31:0] registers_10; // @[Reg_file.scala 20:28]
  reg [31:0] registers_11; // @[Reg_file.scala 20:28]
  reg [31:0] registers_12; // @[Reg_file.scala 20:28]
  reg [31:0] registers_13; // @[Reg_file.scala 20:28]
  reg [31:0] registers_14; // @[Reg_file.scala 20:28]
  reg [31:0] registers_15; // @[Reg_file.scala 20:28]
  reg [31:0] registers_16; // @[Reg_file.scala 20:28]
  reg [31:0] registers_17; // @[Reg_file.scala 20:28]
  reg [31:0] registers_18; // @[Reg_file.scala 20:28]
  reg [31:0] registers_19; // @[Reg_file.scala 20:28]
  reg [31:0] registers_20; // @[Reg_file.scala 20:28]
  reg [31:0] registers_21; // @[Reg_file.scala 20:28]
  reg [31:0] registers_22; // @[Reg_file.scala 20:28]
  reg [31:0] registers_23; // @[Reg_file.scala 20:28]
  reg [31:0] registers_24; // @[Reg_file.scala 20:28]
  reg [31:0] registers_25; // @[Reg_file.scala 20:28]
  reg [31:0] registers_26; // @[Reg_file.scala 20:28]
  reg [31:0] registers_27; // @[Reg_file.scala 20:28]
  reg [31:0] registers_28; // @[Reg_file.scala 20:28]
  reg [31:0] registers_29; // @[Reg_file.scala 20:28]
  wire [31:0] _GEN_1 = 5'h1 == io_r1_addr ? registers_1 : registers_0; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_2 = 5'h2 == io_r1_addr ? registers_2 : _GEN_1; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_3 = 5'h3 == io_r1_addr ? registers_3 : _GEN_2; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_4 = 5'h4 == io_r1_addr ? registers_4 : _GEN_3; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_5 = 5'h5 == io_r1_addr ? registers_5 : _GEN_4; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_6 = 5'h6 == io_r1_addr ? registers_6 : _GEN_5; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_7 = 5'h7 == io_r1_addr ? registers_7 : _GEN_6; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_8 = 5'h8 == io_r1_addr ? registers_8 : _GEN_7; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_9 = 5'h9 == io_r1_addr ? registers_9 : _GEN_8; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_10 = 5'ha == io_r1_addr ? registers_10 : _GEN_9; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_11 = 5'hb == io_r1_addr ? registers_11 : _GEN_10; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_12 = 5'hc == io_r1_addr ? registers_12 : _GEN_11; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_13 = 5'hd == io_r1_addr ? registers_13 : _GEN_12; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_14 = 5'he == io_r1_addr ? registers_14 : _GEN_13; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_15 = 5'hf == io_r1_addr ? registers_15 : _GEN_14; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_16 = 5'h10 == io_r1_addr ? registers_16 : _GEN_15; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_17 = 5'h11 == io_r1_addr ? registers_17 : _GEN_16; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_18 = 5'h12 == io_r1_addr ? registers_18 : _GEN_17; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_19 = 5'h13 == io_r1_addr ? registers_19 : _GEN_18; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_20 = 5'h14 == io_r1_addr ? registers_20 : _GEN_19; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_21 = 5'h15 == io_r1_addr ? registers_21 : _GEN_20; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_22 = 5'h16 == io_r1_addr ? registers_22 : _GEN_21; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_23 = 5'h17 == io_r1_addr ? registers_23 : _GEN_22; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_24 = 5'h18 == io_r1_addr ? registers_24 : _GEN_23; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_25 = 5'h19 == io_r1_addr ? registers_25 : _GEN_24; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_26 = 5'h1a == io_r1_addr ? registers_26 : _GEN_25; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_27 = 5'h1b == io_r1_addr ? registers_27 : _GEN_26; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_28 = 5'h1c == io_r1_addr ? registers_28 : _GEN_27; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  wire [31:0] _GEN_31 = 5'h1 == io_r2_addr ? registers_1 : registers_0; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_32 = 5'h2 == io_r2_addr ? registers_2 : _GEN_31; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_33 = 5'h3 == io_r2_addr ? registers_3 : _GEN_32; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_34 = 5'h4 == io_r2_addr ? registers_4 : _GEN_33; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_35 = 5'h5 == io_r2_addr ? registers_5 : _GEN_34; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_36 = 5'h6 == io_r2_addr ? registers_6 : _GEN_35; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_37 = 5'h7 == io_r2_addr ? registers_7 : _GEN_36; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_38 = 5'h8 == io_r2_addr ? registers_8 : _GEN_37; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_39 = 5'h9 == io_r2_addr ? registers_9 : _GEN_38; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_40 = 5'ha == io_r2_addr ? registers_10 : _GEN_39; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_41 = 5'hb == io_r2_addr ? registers_11 : _GEN_40; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_42 = 5'hc == io_r2_addr ? registers_12 : _GEN_41; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_43 = 5'hd == io_r2_addr ? registers_13 : _GEN_42; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_44 = 5'he == io_r2_addr ? registers_14 : _GEN_43; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_45 = 5'hf == io_r2_addr ? registers_15 : _GEN_44; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_46 = 5'h10 == io_r2_addr ? registers_16 : _GEN_45; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_47 = 5'h11 == io_r2_addr ? registers_17 : _GEN_46; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_48 = 5'h12 == io_r2_addr ? registers_18 : _GEN_47; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_49 = 5'h13 == io_r2_addr ? registers_19 : _GEN_48; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_50 = 5'h14 == io_r2_addr ? registers_20 : _GEN_49; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_51 = 5'h15 == io_r2_addr ? registers_21 : _GEN_50; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_52 = 5'h16 == io_r2_addr ? registers_22 : _GEN_51; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_53 = 5'h17 == io_r2_addr ? registers_23 : _GEN_52; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_54 = 5'h18 == io_r2_addr ? registers_24 : _GEN_53; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_55 = 5'h19 == io_r2_addr ? registers_25 : _GEN_54; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_56 = 5'h1a == io_r2_addr ? registers_26 : _GEN_55; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_57 = 5'h1b == io_r2_addr ? registers_27 : _GEN_56; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  wire [31:0] _GEN_58 = 5'h1c == io_r2_addr ? registers_28 : _GEN_57; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  assign io_r1_data = 5'h1d == io_r1_addr ? registers_29 : _GEN_28; // @[Reg_file.scala 22:20 Reg_file.scala 22:20]
  assign io_r2_data = 5'h1d == io_r2_addr ? registers_29 : _GEN_58; // @[Reg_file.scala 23:20 Reg_file.scala 23:20]
  always @(posedge clock) begin
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h0 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_0 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h1 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_1 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h2 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_2 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h3 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_3 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h4 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_4 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h5 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_5 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h6 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_6 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h7 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_7 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h8 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_8 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h9 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_9 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'ha == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_10 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'hb == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_11 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'hc == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_12 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'hd == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_13 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'he == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_14 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'hf == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_15 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h10 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_16 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h11 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_17 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h12 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_18 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h13 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_19 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h14 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_20 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h15 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_21 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h16 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_22 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h17 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_23 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h18 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_24 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h19 == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_25 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h1a == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_26 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h1b == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_27 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h1c == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_28 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
    if (io_w_en) begin // @[Reg_file.scala 24:22]
      if (5'h1d == io_w_addr) begin // @[Reg_file.scala 25:38]
        registers_29 <= io_w_data; // @[Reg_file.scala 25:38]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  registers_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  registers_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  registers_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  registers_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  registers_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  registers_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  registers_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  registers_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  registers_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  registers_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  registers_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  registers_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  registers_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  registers_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  registers_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  registers_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  registers_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  registers_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  registers_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  registers_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  registers_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  registers_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  registers_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  registers_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  registers_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  registers_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  registers_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  registers_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  registers_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  registers_29 = _RAND_29[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
